module mem_stage (
    input CLK
);
    // 元の riscv_full.v はデータメモリ未実装のため、ここでは何もしません。
endmodule